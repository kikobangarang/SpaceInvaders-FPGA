library ieee;
use ieee.std_logic_1164.all;

entity OutputRegister is
port(	
	D : in std_logic_vector(3 downto 0);
	clk : in std_logic;
	E : in std_logic;
	Reset : in std_logic;
	Q : out std_logic_vector(3 downto 0)
);
end OutputRegister;

architecture behavioral of OutputRegister is

component OutputRegister_FFD port(	
		clk : in std_logic;
		Reset : in std_logic;
		Set : in std_logic;
		D : in std_logic;
		EN : in std_logic;
		Q : out std_logic
);
end component;

begin

FFD_U0: OutputRegister_FFD port map(
		clk => clk,
		Reset => Reset,
		Set => '0',
		D => D(3),
		EN => E,
		Q => Q(3)
);

FFD_U1: OutputRegister_FFD port map(
		clk => clk,
		Reset => Reset,
		Set => '0',
		D => D(2),
		EN => E,
		Q => Q(2)
);

FFD_U2: OutputRegister_FFD port map(
		clk => clk,
		Reset => Reset,
		Set => '0',
		D => D(1),
		EN => E,
		Q => Q(1)
);

FFD_U3: OutputRegister_FFD port map(
		clk => clk,
		Reset => Reset,
		Set => '0',
		D => D(0),
		EN => E,
		Q => Q(0)
);

end behavioral;